library verilog;
use verilog.vl_types.all;
entity t_latch_tb is
end t_latch_tb;
